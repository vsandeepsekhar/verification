`ifndef RAM_SCOREBOARD_SV
`define RAM_SCOREBOARD_SV

class ram_scoreboard extends uvm_scoreboard;

endclass


`endif
