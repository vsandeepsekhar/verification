//--------------------------------------------------------------------------
//This file contains ram config, ram_agent and ram_env class components
//--------------------------------------------------------------------------

`ifdef RAM_AGENT_ENV_CFG__SV
`define RAM_AGENT_ENV_CFG__SV





`endif
